library ieee;
use ieee.std_logic_1164.all;
entity dataPath2 is 
port
(
	
	sel: in std_logic_vector(1 downto 0);
	salida: out std_logic_vector(7 downto 0)
	
);
end dataPath2;

architecture case_arch of dataPath2 is
begin
	process(sel)
	begin
		case (sel) is
			when "00" =>
				salida <= "00000010";
			when "01" =>
				salida <= "00000011";
			when "10" =>
				salida <= "00000100";
			when others =>
				salida <= "00000101";
		end case;
	end process;
end case_arch;


